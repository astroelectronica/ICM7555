.title KiCad schematic
.include "C:/AE/ICM7555/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/ICM7555/_models/C2012X7R2E103K125AA_p.mod"
.include "C:/AE/ICM7555/_models/ICM7555.lib"
R1 /DISC VDD {RDISC}
XU1 0 /TRIGG /OUT VDD /CTRL /TRIGG /DISC VDD ICM7555
R3 /OUT 0 {RLOAD}
R2 /DISC /TRIGG {RTRIGG}
C1 /TRIGG 0 {CTRIGG}
XU3 VDD 0 C2012X7R2A104K125AA_p
V1 VDD 0 {VSUPPLY}
XU2 /CTRL 0 C2012X7R2E103K125AA_p
.end
